`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: _5WB
// Description: 
//////////////////////////////////////////////////////////////////////////////////


module _5WB(

    );
endmodule
