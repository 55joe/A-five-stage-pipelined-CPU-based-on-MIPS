module _0InstructionMemory(
	input      [32 -1:0] Address, 
	output reg [32 -1:0] Instruction
);
	
	initial
		Instruction = 32'b0;

	always @(*)
		case (Address[10:2])
/*
9'd0:  Instruction <= 32'b00100000000111010000001000000000;
9'd1:  Instruction <= 32'b00100000000100000000000000000001;
9'd2:  Instruction <= 32'b10001100000001010000000000000000;
9'd3:  Instruction <= 32'b00100000000001000000000000000100;
9'd4:  Instruction <= 32'b00001100000100000000000001000010;
9'd5:  Instruction <= 32'b00000000000000000000000000000000;
9'd6:  Instruction <= 32'b00001000000100000000000001010011;
9'd7:  Instruction <= 32'b00000000000000000000000000000000;
9'd8:  Instruction <= 32'b00100000000000010000000000000100;
9'd9:  Instruction <= 32'b00000011101000011110100000100010;
9'd10: Instruction <= 32'b10101111101111110000000000000000;
9'd11: Instruction <= 32'b00000001000000000100100000100000;
9'd12: Instruction <= 32'b00100000000000010000000000000001;
9'd13: Instruction <= 32'b00000001001000010100100000100010;
9'd14: Instruction <= 32'b00000001000000000101000000100000;
9'd15: Instruction <= 32'b00000000000010100101000010000000;
9'd16: Instruction <= 32'b00000000100010101100000000100000;
9'd17: Instruction <= 32'b10001111000010110000000000000000;
9'd18: Instruction <= 32'b00100010000100000000000000000001;
9'd19: Instruction <= 32'b00000001001000000101000000100000;
9'd20: Instruction <= 32'b00000000000010100101000010000000;
9'd21: Instruction <= 32'b00000000100010101100000000100000;
9'd22: Instruction <= 32'b10001111000011000000000000000000;
9'd23: Instruction <= 32'b00000001011011000000100000101010;
9'd24: Instruction <= 32'b00010000001000000000000000000111;
9'd25: Instruction <= 32'b00000000000000000000000000000000;
9'd26: Instruction <= 32'b00100000000000010000000000000001;
9'd27: Instruction <= 32'b00000001001000010100100000100010;
9'd28: Instruction <= 32'b00000101001000000000000000000011;
9'd29: Instruction <= 32'b00000000000000000000000000000000;
9'd30: Instruction <= 32'b00001000000100000000000000010010;
9'd31: Instruction <= 32'b00000000000000000000000000000000;
9'd32: Instruction <= 32'b00100001001000100000000000000001;
9'd33: Instruction <= 32'b10001111101111110000000000000000;
9'd34: Instruction <= 32'b00100011101111010000000000000100;
9'd35: Instruction <= 32'b00000011111000000000000000001000;
9'd36: Instruction <= 32'b00000000000000000000000000000000;
9'd37: Instruction <= 32'b00100000000000010000000000000100;
9'd38: Instruction <= 32'b00000011101000011110100000100010;
9'd39: Instruction <= 32'b10101111101111110000000000000000;
9'd40: Instruction <= 32'b00000001000000000110100000100000;
9'd41: Instruction <= 32'b00100000000000010000000000000001;
9'd42: Instruction <= 32'b00000001101000010110100000100010;
9'd43: Instruction <= 32'b00000001000000000111000000100000;
9'd44: Instruction <= 32'b00000000000010000111000010000000;
9'd45: Instruction <= 32'b00000000100011100100100000100000;
9'd46: Instruction <= 32'b10001101001011110000000000000000;
9'd47: Instruction <= 32'b00000001101000001100100000100000;
9'd48: Instruction <= 32'b00000000000110011100100010000000;
9'd49: Instruction <= 32'b00100011001110000000000000000100;
9'd50: Instruction <= 32'b00000000100110000100100000100000;
9'd51: Instruction <= 32'b00000000100110010101000000100000;
9'd52: Instruction <= 32'b10001101010010110000000000000000;
9'd53: Instruction <= 32'b10101101001010110000000000000000;
9'd54: Instruction <= 32'b00100000000000010000000000000001;
9'd55: Instruction <= 32'b00000001101000010110100000100010;
9'd56: Instruction <= 32'b00000001101001100000100000101010;
9'd57: Instruction <= 32'b00010000001000001111111111110101;
9'd58: Instruction <= 32'b00000000000000000000000000000000;
9'd59: Instruction <= 32'b00000000000001100011000010000000;
9'd60: Instruction <= 32'b00000000100001100100100000100000;
9'd61: Instruction <= 32'b10101101001011110000000000000000;
9'd62: Instruction <= 32'b10001111101111110000000000000000;
9'd63: Instruction <= 32'b00100011101111010000000000000100;
9'd64: Instruction <= 32'b00000011111000000000000000001000;
9'd65: Instruction <= 32'b00000000000000000000000000000000;
9'd66: Instruction <= 32'b00100000000000010000000000000100;
9'd67: Instruction <= 32'b00000011101000011110100000100010;
9'd68: Instruction <= 32'b10101111101111110000000000000000;
9'd69: Instruction <= 32'b00100000000010000000000000000001;
9'd70: Instruction <= 32'b00001100000100000000000000001000;
9'd71: Instruction <= 32'b00000000000000000000000000000000;
9'd72: Instruction <= 32'b00000000010000000011000000100000;
9'd73: Instruction <= 32'b00001100000100000000000000100101;
9'd74: Instruction <= 32'b00000000000000000000000000000000;
9'd75: Instruction <= 32'b00100001000010000000000000000001;
9'd76: Instruction <= 32'b00000001000001010000100000101010;
9'd77: Instruction <= 32'b00010100001000001111111111111000;
9'd78: Instruction <= 32'b00000000000000000000000000000000;
9'd79: Instruction <= 32'b10001111101111110000000000000000;
9'd80: Instruction <= 32'b00100011101111010000000000000100;
9'd81: Instruction <= 32'b00000011111000000000000000001000;
9'd82: Instruction <= 32'b00000000000000000000000000000000;
9'd83: Instruction <= 32'b00000000000000000000000000000000;
*/
9'd0: Instruction <= 32'h201d0200;
9'd1: Instruction <= 32'h20100001;
9'd2: Instruction <= 32'h8c050000;
9'd3: Instruction <= 32'h20040004;
9'd4: Instruction <= 32'h0c100042;
9'd5: Instruction <= 32'h00000000;
9'd6: Instruction <= 32'h08100053;
9'd7: Instruction <= 32'h00000000;
9'd8: Instruction <= 32'h20010004;
9'd9: Instruction <= 32'h03a1e822;
9'd10: Instruction <= 32'hafbf0000;
9'd11: Instruction <= 32'h01004820;
9'd12: Instruction <= 32'h20010001;
9'd13: Instruction <= 32'h01214822;
9'd14: Instruction <= 32'h01005020;
9'd15: Instruction <= 32'h000a5080;
9'd16: Instruction <= 32'h008ac020;
9'd17: Instruction <= 32'h8f0b0000;
9'd18: Instruction <= 32'h22100001;
9'd19: Instruction <= 32'h01205020;
9'd20: Instruction <= 32'h000a5080;
9'd21: Instruction <= 32'h008ac020;
9'd22: Instruction <= 32'h8f0c0000;
9'd23: Instruction <= 32'h016c082a;
9'd24: Instruction <= 32'h10200007;
9'd25: Instruction <= 32'h00000000;
9'd26: Instruction <= 32'h20010001;
9'd27: Instruction <= 32'h01214822;
9'd28: Instruction <= 32'h05200003;
9'd29: Instruction <= 32'h00000000;
9'd30: Instruction <= 32'h08100012;
9'd31: Instruction <= 32'h00000000;
9'd32: Instruction <= 32'h21220001;
9'd33: Instruction <= 32'h8fbf0000;
9'd34: Instruction <= 32'h23bd0004;
9'd35: Instruction <= 32'h03e00008;
9'd36: Instruction <= 32'h00000000;
9'd37: Instruction <= 32'h20010004;
9'd38: Instruction <= 32'h03a1e822;
9'd39: Instruction <= 32'hafbf0000;
9'd40: Instruction <= 32'h01006820;
9'd41: Instruction <= 32'h20010001;
9'd42: Instruction <= 32'h01a16822;
9'd43: Instruction <= 32'h01007020;
9'd44: Instruction <= 32'h00087080;
9'd45: Instruction <= 32'h008e4820;
9'd46: Instruction <= 32'h8d2f0000;
9'd47: Instruction <= 32'h01a0c820;
9'd48: Instruction <= 32'h0019c880;
9'd49: Instruction <= 32'h23380004;
9'd50: Instruction <= 32'h00984820;
9'd51: Instruction <= 32'h00995020;
9'd52: Instruction <= 32'h8d4b0000;
9'd53: Instruction <= 32'had2b0000;
9'd54: Instruction <= 32'h20010001;
9'd55: Instruction <= 32'h01a16822;
9'd56: Instruction <= 32'h01a6082a;
9'd57: Instruction <= 32'h1020fff5;
9'd58: Instruction <= 32'h00000000;
9'd59: Instruction <= 32'h00063080;
9'd60: Instruction <= 32'h00864820;
9'd61: Instruction <= 32'had2f0000;
9'd62: Instruction <= 32'h8fbf0000;
9'd63: Instruction <= 32'h23bd0004;
9'd64: Instruction <= 32'h03e00008;
9'd65: Instruction <= 32'h00000000;
9'd66: Instruction <= 32'h20010004;
9'd67: Instruction <= 32'h03a1e822;
9'd68: Instruction <= 32'hafbf0000;
9'd69: Instruction <= 32'h20080001;
9'd70: Instruction <= 32'h0c100008;
9'd71: Instruction <= 32'h00000000;
9'd72: Instruction <= 32'h00403020;
9'd73: Instruction <= 32'h0c100025;
9'd74: Instruction <= 32'h00000000;
9'd75: Instruction <= 32'h21080001;
9'd76: Instruction <= 32'h0105082a;
9'd77: Instruction <= 32'h1420fff8;
9'd78: Instruction <= 32'h00000000;
9'd79: Instruction <= 32'h8fbf0000;
9'd80: Instruction <= 32'h23bd0004;
9'd81: Instruction <= 32'h03e00008;
9'd82: Instruction <= 32'h00000000;
9'd83: Instruction <= 32'h00000000;
9'd84: Instruction <= 32'h8c040000;
9'd85: Instruction <= 32'h20840001;
9'd86: Instruction <= 32'h3c054000;
9'd87: Instruction <= 32'h20a50010;
9'd88: Instruction <= 32'h200603e8;
9'd89: Instruction <= 32'h20071f40;
9'd90: Instruction <= 32'h20080000;
9'd91: Instruction <= 32'h21080001;
9'd92: Instruction <= 32'h1104fff6;
9'd93: Instruction <= 32'h00000000;
9'd94: Instruction <= 32'h00084080;
9'd95: Instruction <= 32'h8d090000;
9'd96: Instruction <= 32'h00084082;
9'd97: Instruction <= 32'h200a0000;
9'd98: Instruction <= 32'haca90000;
9'd99: Instruction <= 32'h214a0001;
9'd100: Instruction <= 32'h1147fff6;
9'd101: Instruction <= 32'h00000000;
9'd102: Instruction <= 32'h200b0000;
9'd103: Instruction <= 32'h216b0001;
9'd104: Instruction <= 32'h1566fffe;
9'd105: Instruction <= 32'h00000000;
9'd106: Instruction <= 32'h20170001;
9'd107: Instruction <= 32'h00176880;
9'd108: Instruction <= 32'h01a56820;
9'd109: Instruction <= 32'h8dae0000;
9'd110: Instruction <= 32'h0c100091;
9'd111: Instruction <= 32'h00000000;
9'd112: Instruction <= 32'h200b0000;
9'd113: Instruction <= 32'h216b0001;
9'd114: Instruction <= 32'h1566fffe;
9'd115: Instruction <= 32'h00000000;
9'd116: Instruction <= 32'h20170002;
9'd117: Instruction <= 32'h00176880;
9'd118: Instruction <= 32'h01a56820;
9'd119: Instruction <= 32'h8dae0000;
9'd120: Instruction <= 32'h0c100091;
9'd121: Instruction <= 32'h00000000;
9'd122: Instruction <= 32'h200b0000;
9'd123: Instruction <= 32'h216b0001;
9'd124: Instruction <= 32'h1566fffe;
9'd125: Instruction <= 32'h00000000;
9'd126: Instruction <= 32'h20170003;
9'd127: Instruction <= 32'h00176880;
9'd128: Instruction <= 32'h01a56820;
9'd129: Instruction <= 32'h8dae0000;
9'd130: Instruction <= 32'h0c100091;
9'd131: Instruction <= 32'h00000000;
9'd132: Instruction <= 32'h200b0000;
9'd133: Instruction <= 32'h216b0001;
9'd134: Instruction <= 32'h1566fffe;
9'd135: Instruction <= 32'h00000000;
9'd136: Instruction <= 32'h20170004;
9'd137: Instruction <= 32'h00176880;
9'd138: Instruction <= 32'h01a56820;
9'd139: Instruction <= 32'h8dae0000;
9'd140: Instruction <= 32'h0c100091;
9'd141: Instruction <= 32'h00000000;
9'd142: Instruction <= 32'h200b0000;
9'd143: Instruction <= 32'h08100063;
9'd144: Instruction <= 32'h00000000;
9'd145: Instruction <= 32'h20010004;
9'd146: Instruction <= 32'h03a1e822;
9'd147: Instruction <= 32'hafbf0000;
9'd148: Instruction <= 32'h15c0000a;
9'd149: Instruction <= 32'h00000000;
9'd150: Instruction <= 32'h20100001;
9'd151: Instruction <= 32'h20110001;
9'd152: Instruction <= 32'h20120001;
9'd153: Instruction <= 32'h20130001;
9'd154: Instruction <= 32'h20140001;
9'd155: Instruction <= 32'h20150001;
9'd156: Instruction <= 32'h20160000;
9'd157: Instruction <= 32'h0810016b;
9'd158: Instruction <= 32'h00000000;
9'd159: Instruction <= 32'h20010001;
9'd160: Instruction <= 32'h01c17022;
9'd161: Instruction <= 32'h15c0000a;
9'd162: Instruction <= 32'h00000000;
9'd163: Instruction <= 32'h20100000;
9'd164: Instruction <= 32'h20110001;
9'd165: Instruction <= 32'h20120001;
9'd166: Instruction <= 32'h20130000;
9'd167: Instruction <= 32'h20140000;
9'd168: Instruction <= 32'h20150000;
9'd169: Instruction <= 32'h20160000;
9'd170: Instruction <= 32'h0810016b;
9'd171: Instruction <= 32'h00000000;
9'd172: Instruction <= 32'h20010001;
9'd173: Instruction <= 32'h01c17022;
9'd174: Instruction <= 32'h15c0000a;
9'd175: Instruction <= 32'h00000000;
9'd176: Instruction <= 32'h20100001;
9'd177: Instruction <= 32'h20110001;
9'd178: Instruction <= 32'h20120000;
9'd179: Instruction <= 32'h20130001;
9'd180: Instruction <= 32'h20140001;
9'd181: Instruction <= 32'h20150000;
9'd182: Instruction <= 32'h20160001;
9'd183: Instruction <= 32'h0810016b;
9'd184: Instruction <= 32'h00000000;
9'd185: Instruction <= 32'h20010001;
9'd186: Instruction <= 32'h01c17022;
9'd187: Instruction <= 32'h15c0000a;
9'd188: Instruction <= 32'h00000000;
9'd189: Instruction <= 32'h20100001;
9'd190: Instruction <= 32'h20110001;
9'd191: Instruction <= 32'h20120001;
9'd192: Instruction <= 32'h20130001;
9'd193: Instruction <= 32'h20140000;
9'd194: Instruction <= 32'h20150000;
9'd195: Instruction <= 32'h20160001;
9'd196: Instruction <= 32'h0810016b;
9'd197: Instruction <= 32'h00000000;
9'd198: Instruction <= 32'h20010001;
9'd199: Instruction <= 32'h01c17022;
9'd200: Instruction <= 32'h15c0000a;
9'd201: Instruction <= 32'h00000000;
9'd202: Instruction <= 32'h20100000;
9'd203: Instruction <= 32'h20110001;
9'd204: Instruction <= 32'h20120001;
9'd205: Instruction <= 32'h20130000;
9'd206: Instruction <= 32'h20140000;
9'd207: Instruction <= 32'h20150001;
9'd208: Instruction <= 32'h20160001;
9'd209: Instruction <= 32'h0810016b;
9'd210: Instruction <= 32'h00000000;
9'd211: Instruction <= 32'h20010001;
9'd212: Instruction <= 32'h01c17022;
9'd213: Instruction <= 32'h15c0000a;
9'd214: Instruction <= 32'h00000000;
9'd215: Instruction <= 32'h20100001;
9'd216: Instruction <= 32'h20110000;
9'd217: Instruction <= 32'h20120001;
9'd218: Instruction <= 32'h20130001;
9'd219: Instruction <= 32'h20140000;
9'd220: Instruction <= 32'h20150001;
9'd221: Instruction <= 32'h20160001;
9'd222: Instruction <= 32'h0810016b;
9'd223: Instruction <= 32'h00000000;
9'd224: Instruction <= 32'h20010001;
9'd225: Instruction <= 32'h01c17022;
9'd226: Instruction <= 32'h15c0000a;
9'd227: Instruction <= 32'h00000000;
9'd228: Instruction <= 32'h20100001;
9'd229: Instruction <= 32'h20110000;
9'd230: Instruction <= 32'h20120001;
9'd231: Instruction <= 32'h20130001;
9'd232: Instruction <= 32'h20140001;
9'd233: Instruction <= 32'h20150001;
9'd234: Instruction <= 32'h20160001;
9'd235: Instruction <= 32'h0810016b;
9'd236: Instruction <= 32'h00000000;
9'd237: Instruction <= 32'h20010001;
9'd238: Instruction <= 32'h01c17022;
9'd239: Instruction <= 32'h15c0000a;
9'd240: Instruction <= 32'h00000000;
9'd241: Instruction <= 32'h20100001;
9'd242: Instruction <= 32'h20110001;
9'd243: Instruction <= 32'h20120001;
9'd244: Instruction <= 32'h20130000;
9'd245: Instruction <= 32'h20140000;
9'd246: Instruction <= 32'h20150000;
9'd247: Instruction <= 32'h20160000;
9'd248: Instruction <= 32'h0810016b;
9'd249: Instruction <= 32'h00000000;
9'd250: Instruction <= 32'h20010001;
9'd251: Instruction <= 32'h01c17022;
9'd252: Instruction <= 32'h15c0000a;
9'd253: Instruction <= 32'h00000000;
9'd254: Instruction <= 32'h20100001;
9'd255: Instruction <= 32'h20110001;
9'd256: Instruction <= 32'h20120001;
9'd257: Instruction <= 32'h20130001;
9'd258: Instruction <= 32'h20140001;
9'd259: Instruction <= 32'h20150001;
9'd260: Instruction <= 32'h20160001;
9'd261: Instruction <= 32'h0810016b;
9'd262: Instruction <= 32'h00000000;
9'd263: Instruction <= 32'h20010001;
9'd264: Instruction <= 32'h01c17022;
9'd265: Instruction <= 32'h15c0000a;
9'd266: Instruction <= 32'h00000000;
9'd267: Instruction <= 32'h20100001;
9'd268: Instruction <= 32'h20110001;
9'd269: Instruction <= 32'h20120001;
9'd270: Instruction <= 32'h20130001;
9'd271: Instruction <= 32'h20140000;
9'd272: Instruction <= 32'h20150001;
9'd273: Instruction <= 32'h20160001;
9'd274: Instruction <= 32'h0810016b;
9'd275: Instruction <= 32'h00000000;
9'd276: Instruction <= 32'h20010001;
9'd277: Instruction <= 32'h01c17022;
9'd278: Instruction <= 32'h15c0000a;
9'd279: Instruction <= 32'h00000000;
9'd280: Instruction <= 32'h20100001;
9'd281: Instruction <= 32'h20110001;
9'd282: Instruction <= 32'h20120001;
9'd283: Instruction <= 32'h20130000;
9'd284: Instruction <= 32'h20140001;
9'd285: Instruction <= 32'h20150001;
9'd286: Instruction <= 32'h20160001;
9'd287: Instruction <= 32'h0810016b;
9'd288: Instruction <= 32'h00000000;
9'd289: Instruction <= 32'h20010001;
9'd290: Instruction <= 32'h01c17022;
9'd291: Instruction <= 32'h15c0000a;
9'd292: Instruction <= 32'h00000000;
9'd293: Instruction <= 32'h20100000;
9'd294: Instruction <= 32'h20110000;
9'd295: Instruction <= 32'h20120001;
9'd296: Instruction <= 32'h20130001;
9'd297: Instruction <= 32'h20140001;
9'd298: Instruction <= 32'h20150001;
9'd299: Instruction <= 32'h20160001;
9'd300: Instruction <= 32'h0810016b;
9'd301: Instruction <= 32'h00000000;
9'd302: Instruction <= 32'h20010001;
9'd303: Instruction <= 32'h01c17022;
9'd304: Instruction <= 32'h15c0000a;
9'd305: Instruction <= 32'h00000000;
9'd306: Instruction <= 32'h20100001;
9'd307: Instruction <= 32'h20110000;
9'd308: Instruction <= 32'h20120000;
9'd309: Instruction <= 32'h20130001;
9'd310: Instruction <= 32'h20140001;
9'd311: Instruction <= 32'h20150001;
9'd312: Instruction <= 32'h20160000;
9'd313: Instruction <= 32'h0810016b;
9'd314: Instruction <= 32'h00000000;
9'd315: Instruction <= 32'h20010001;
9'd316: Instruction <= 32'h01c17022;
9'd317: Instruction <= 32'h15c0000a;
9'd318: Instruction <= 32'h00000000;
9'd319: Instruction <= 32'h20100000;
9'd320: Instruction <= 32'h20110001;
9'd321: Instruction <= 32'h20120001;
9'd322: Instruction <= 32'h20130001;
9'd323: Instruction <= 32'h20140001;
9'd324: Instruction <= 32'h20150000;
9'd325: Instruction <= 32'h20160001;
9'd326: Instruction <= 32'h0810016b;
9'd327: Instruction <= 32'h00000000;
9'd328: Instruction <= 32'h20010001;
9'd329: Instruction <= 32'h01c17022;
9'd330: Instruction <= 32'h15c0000a;
9'd331: Instruction <= 32'h00000000;
9'd332: Instruction <= 32'h20100001;
9'd333: Instruction <= 32'h20110000;
9'd334: Instruction <= 32'h20120000;
9'd335: Instruction <= 32'h20130001;
9'd336: Instruction <= 32'h20140001;
9'd337: Instruction <= 32'h20150001;
9'd338: Instruction <= 32'h20160001;
9'd339: Instruction <= 32'h0810016b;
9'd340: Instruction <= 32'h00000000;
9'd341: Instruction <= 32'h20010001;
9'd342: Instruction <= 32'h01c17022;
9'd343: Instruction <= 32'h15c0000c;
9'd344: Instruction <= 32'h00000000;
9'd345: Instruction <= 32'h20010001;
9'd346: Instruction <= 32'h01c17022;
9'd347: Instruction <= 32'h20100001;
9'd348: Instruction <= 32'h20110000;
9'd349: Instruction <= 32'h20120000;
9'd350: Instruction <= 32'h20130000;
9'd351: Instruction <= 32'h20140001;
9'd352: Instruction <= 32'h20150001;
9'd353: Instruction <= 32'h20160001;
9'd354: Instruction <= 32'h0810016b;
9'd355: Instruction <= 32'h00000000;
9'd356: Instruction <= 32'h20100000;
9'd357: Instruction <= 32'h20110000;
9'd358: Instruction <= 32'h20120000;
9'd359: Instruction <= 32'h20130000;
9'd360: Instruction <= 32'h20140000;
9'd361: Instruction <= 32'h20150000;
9'd362: Instruction <= 32'h20160000;
9'd363: Instruction <= 32'h8fbf0000;
9'd364: Instruction <= 32'h23bd0004;
9'd365: Instruction <= 32'h03e00008;
9'd366: Instruction <= 32'h00000000;




default:Instruction <= 32'b0;


		endcase
		
endmodule
