`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: _stall
// Description:
//////////////////////////////////////////////////////////////////////////////////


module _stall(
    input wire clk,
    input wire rst,
    input wire stall_load,
    output wire stall
    );

assign stall = stall_load;


endmodule
